module CTRL_weight_reload #(
    parameters
) (
    input wire we_rl,
    output wire 
);
    
endmodule